module first_project
(
input in,
output out
);

assign out = in
endmodule;